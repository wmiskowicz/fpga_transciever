interface rx_in_if ();
  logic               clk;
  logic         [7:0] rxd;
  logic               rxdv;
  logic               rxer;
endinterface
